`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DtbuQpcJqp26T+zectVGkmv5OK4mWShIpEVedtenQO4zrfts4wM74T3k9nKrxxt2W1tPWM0Wmnk1
Z8OCLhrM3g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d2i3th88eOgh94cMcBowDLISEdIQpnbxArCBVrpPX/HD4Zgsxjhba3lHOSbEcBQEOXI1mqJjQscR
sBrCpTdJP4j+/6ewEaQd7mINh2Z8/E3qYQ1sA3rw/B8unw8l+smmrHSMjvkG0HESDch2UYD6DiOd
DnzkOUhdr306BpIEWzA=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ILjvPSvbnKoV5EUyxxfwvyzjsMxc+lZdcOt0ULYWf2ZmnkElI+JyAfmZ566Cv5BybvIAbpkE4TAs
lbFdJpKI0wxt0RVWOuWLyVmxuNoSdo4QruYKvQVHEs1XVTIuysBzqE/vE45srqQBFh0chx3HuYsH
25NRSNvvSDfGVSbPt2Y=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DJLt4ZDDim1Hm/RC/uN3S28HGocmb+fp1NEHpBa1fctdY6Xa0dl9swUDB43bBqke6rH6S+aVFKvY
+VIXG+GN10oOrqBtTUlx2bph1/JtHXfdxrD/iDoM9kZAd44aYFcDDXx5Sf/dv44DWtk6Y6F1mpl8
JLJskCz/HtLXPFpjgPBR2FayX3lU5het3dp8+v5TVMXYmTNhbfbjiZapWjulNJHmNNgQh/0OXg9g
CVaGlzLERyylDYSPUDRiEjaCHzGk4TJIFiaR22AQL3bMyQcJgf9vV+5cq/llII6IkC1zQQzMnX0F
zMKS9e70V56XKvWAZvl54nsh7HNf4hYe1RK93w==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dFBNohZIkCMhAoWOoktwYbWbF2tqJ762dUmpci7xJH+4DC2zZzFfQHC8adbAxdiNfNknj7dcVe2+
kEiX/hxC5LNOFwVUPriXwk4eC/0JE9Q0cKzIC42UDbXN7Gh+mUzPwxacEVqKG6pxmwgmw54Y+3qw
tPeM0v0WWchQeXuu8sLzfhAHySx759Rnmac039Bizpezjo6EzBHljszn7OSgYTMFlkPkF/xWBRbr
PtbvLsmJ77wKiJgiwrzsx00eSzHRPntQzHpul8zDvJ7GWVDjDYs1KxV+W+K5EbdA+VhVXdTfalgE
da0UFM277buLz6cWMHPipRcZ1BQpXoyLfH0Ntg==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M7cBjZ4oaFyC5MJnXQ2hoTYtu56oRbTi39VhEd3XwNgykupeLNWKfnTaF1F5XjkTEK+u7OKGP9b+
BPwvCCeyRMGToU3e6f+038OgCktGUmYR5K8IOq6/L1wdzi0fvinc2ZcnXygxPvS9CwChP6kQ+3nA
z3lVzCic6EARe4sKkUYVCLiIsTNc36CDJJnh3n7GyYLy7bhkSP481skgtiNmP7z/q+dfYYSqocgG
yETWD5QhiI2jRRuc3W3herl668378xA/1BlvNKK69Jlnh2n0iQg6i/b2AvKdgoCN0zpAv462oTKA
BO8Lpw0sSopNxXj/MEgPTpC3/+fRT4TdCtIYLA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5824)
`protect data_block
TkXIcuaIIkxkfSuRsCApwrY4vCIjc00cl+AeozJME8Kx8ueNQHDxoUpcFiDj9gSELrLE1VaWVz8b
mveGHs3Aa6ZzcT+diZh2qZfMSQ98atsFREfgTwykuu68SCX8IAv0Xz1t1R+Otn/BZey+OaeZl/YC
pNh44zEDeg9s2TfTr/sWqkBCOs1/nAeF03BpXqQytT38yWMH502VUCAfCR0I3j9eAGrrJ6tfd6kM
izJPZ38ZpO+iy8kg7iisGIQA7/iHYnTgMsbDu+laXHm592vl/uDzX5lOBfTmt5PiG5hQ3LZ6aUE5
kLnke4Pab2daY8B30banap9KzWlmdNc78zLWYdkZbRKROtsfSGU7uhxxyH2RVjOw0e9sa5shy0ie
uJdBH2Aku204uzZxmO0b3e8YUOTrdys8Hq/keI0zN6d/uKQ32RWney2AxJNr8xNQb68LezbpOQYU
GsY9ZSyKgdTjXNiWdv6wxOZPGLLZpztgej6ZvfP8e/pY5VMWqHspiLzxkd9/TDvQMegnQf8Z80ZT
vbte+cSwmXyS0SXKYBjFG5M0BYmfsuEqqOFgzYn08NWqeoAHAxPhsakEx34/abeHW6krNBRlywBt
UpxSX2uip+vLRCd3nyQECFT+YS9mjcwQkGv4IYFcDosALTt3eMFCT3/1ylWPewM1ku4fV+tvA86q
Dt3gW80+HTijHU0g9+MgkRMuvNW4YhTqldakSQ/h+ce2jOd5tnaCbnRofqX4vpC9eX/I4whBmMZB
zzMz/8c6xfM2Nu7iRwLhBcH8zKjegbKM8LNxGBJZo67DLX9fep/Zz9JJG/6OxiJRx3cP/D0mIkMU
gw67f+263lZPz0A05hG285S44g6aPD0e75VDs+sq07bJ8fuqeU2HGDcoSvyG1y1ry1Ywol3Q5mY2
qdk/jcldvCSqAs8dvL7ZGV6wk5GgjBJGQAz/XVpVdrMYVvYBdGbKijseXdyFRJHX/pkQnQ2GcP+9
PVYK7KwiWvC0SlL63zKdM792YwxuynxFi9zlkSv4r8PzCQKfCTU7IfYNauj2OSOA5izuOZLUlCQa
igapF8FAaC4dIVZcuZly/xDBCPz138LR3KVjqgb9gzLwaOTrgwm7YixHW2Kw+tGGXxIpLZvHkC0P
FEE8BzUqa2WopWrtaE+PZkHMaVWIAlrcy/HVi56FU8x9q469vrB9w/WFDqcO/Ge5KWVpwHrNos8N
TkZeOfsKxs5CvGCytgeCjX8oIz5Zwi53Ka3ni3pD5JmYkXVr2kIJ3uUuXgCvxYGtmmKjzNaTE/p5
fkhVdh7ljETVF/1Tnka0wS2o/0AmzCYMvRPcPxX1HDM6a9FatzyfM2lqszEhZj73UeINJGhiUrGh
ATPz7/2vC0EP5zwrsc6MHDlNn2w5dQsoUSriOQbmWNm0ipXkWE7Wpi5PnIVhKFH2uvWMoof68kfm
56Jx2o0y7vaunFz/nGtKd6x/BLtUXhzdqovupNAUC1h1X9kf9dH600YphcQNGMsMARt/KOBeKqU/
W3iKZOUtw4PG8HEi12OysaehpD0n0Y/+C8MX2xN1fG6w4t/Vhav5ay6iygWl8LpuKkJBsvAyoJyN
jv+713v2qyc9PE4scHdCLGGHYqwnMCDmm/H1ua++zm3s6NYu80OxUjqEdVzwWzS63VoxOkPKaNZs
r1toBY2pQBGs9DX//ToZEnPWKqMI8WahgNdy57cbZtclfBbiLGcXCXneBW5fLKflFmVSAU76TXx+
LG8rVbXTkLPiRhWzriswmyFHU7KqpIIPA2hTDymFCdYFSaGhXC8TXs3p3rWSNMpMfoSfAX6+X0zP
11QY01s5pHesnQLlCE6gK0DmlBgdAwbV/LY/IKfcyWyHdliFLWfdvCOQJxtUwsmx4VCH1wgGEESA
qfbPx4Ixh3tNDQRTHmWgjCA1uG2VkOFuXNywGGwMFtcbQj1b1H1Ql3Jx2JOdijKPUCduliKNCIKu
2kiRNNfC0zXdL67XsV+HQAWuykL9OUw8zxWNBD5Ti2qZp8pQLUKq42/v+1CCOObPdVWBnRpm3CE4
6cUDe823Zq5ANqX8pvf9lw8Qdq3w0B+l+iEqaxNhG7sVQg7WiT9Q2TLU739IvfT4HkU++Z0rvhTX
Rfut5pu1s0tU1K2EuT/7UhTMYVbzelGBt3FZq/SJPy7qS4R3j0wlfYeTd4XAbgYGCrl9vMyNx51y
2jPFx+No7y72jO6VGF5fbTpupoopKdZvTUVed0q7QrwO7NC0s/8Ob29stqKiK6mdpsBZj7f5IRgZ
VdepuF7EsTDcDiVdQAUrAQf9ir3bopnCx+OdR0d5QNPnBkU2bhYFEfKG+EKqS92s0mT2/dE0Rhp7
Xd9NAa+PRyQXOrTWUCGXP532bQv2T1le3SR7CKruV/0rEDAr+qaj/1HIO/LshX4ziB4iSuQZ2HB3
YWxC4fcX4zHnoHMN4H9lXdb7/KBZhOIrH4f4/DtefK8M2UO7fM6bw9b9OT1fKrBKQ3XB1cb3pA3b
2r0Y0IsKpaQauiIemzLfQ2Y/EbhJ38vv/ikgfUnH4puw++yRFqLzCEHnCbuBXG5RHLtNASL3T3yL
wVlldPXbGWKg4S6TDALPNaYPVd4QuPkXiLl4ubD3f0aTeemIsWIBt3AIDJ6GXJ8kcHYNruHMeuRk
DFq/KCUp6xl9rOf1rlzTAcu7Ff8R6sCW38TKMGGmq7ZMdSYfblJUTITk5/seEDHWuIWqyhAdZUJd
X5LNCFhf6v3kemTAZ6B1nW8hHz88X4Zy9D5R6jZvzAZvHgqC67QXJIS8SFMRGF0++JC861T5p5oj
roXbsQn5e9FPgia/re5hYbA3xVuS/f2/il/9ode7Uw8unKZLEj5nJzLIhK2kotAC84dHlc18OcOq
iU8luPRxLyTz0sY5JGUq9Kw7+HYR2EtSEfvV28mm8kQKa7a7bHawfWYi55akpFxUJKmmHVirV1Jl
fLpieSvS0A/o0HywNSME+j3z6ZAyk+AnBq/n/p5zHzP7CnZ7U4mWELJ/ALsYjHt0WA+R64QF+0JE
mhgv1Vxeq6r6fPx0BJ0g3cAeev+6xWQpR6IYnMiTpYzoHEW37yFmqcXNumM072eqSonj9FkGqllk
nswk857z3qbRIPjdHMMnzx+MZmAbteX27NbAShbPGRZpORb/VZ/L3qHqcvHhSHvcr6zWiQR1WLxo
2HoZq9jV1Uv6J4cHWc3TyxEPgn15YBc6r+kIBMQdrgA8gUXXVBuUvnhTiiZei1VP3BygINkXW60g
n/8MayokKRqkB21K+p8WlAT6IJVPFm4+CehrtTgx7iPSN6+4Ix5QEnsjfC211VrISJdpargZRdwf
IIIC1+rniSNhNHcBzuQg6WX1Ps0C/CSrqCdjZ+kEDsj7oMwHLj3T1s2DCcNdMy1RjaS3PBXk5Y//
W4YGAF25ZvXPposSzZt5rdBCcOweTeXPvS1CKxZjc+0itg8JwZ64yrxOyE+/2eLQ5ixZWz/FVN38
nGXmaKWqc+euZ5XrzN4MB46TJJ5/bjPpu5NVHsfE66N/EyrQzuC+sT+1p1a1UF5aNiVNn87MSueS
tZDf9oJCmD3CD9jrGEqqq7EVf8GgruiAnbP1rcTwnaJOll3xrYEF8aVfUyYNWVbjzLOc5/YYtIGv
8LRZ0TxoxcK8IXmdPT0kcD4F6nOl0qpB1vNIk92FUo2SiCNiErmTtb9dB9eSwcWDb3TMAcHhDb61
ugaIFFYG+WLhvEQ2c2BVBWm4jwa/mWbJ9vMIwvhRCTit7mf7n86h76DQsAtipJmPTgmKpURIzhg2
XaWQoik7IbKnyWt94NkqtFenoKFNDFGtWd+m7z+Gx2xc1QiiYm9fHVN8SvPGotNn1KMmBqEAK7oW
yfFX5Xvi1Q21QsA+ALDs8khGMpms5ziZCS3d6y2m0qxexquOIN3NH1e8Hrq8wYsl4TTnqCB3sbTf
PJTrRJAoDgfKlPu0WTcEd95GYEbUGElJLlPrnZ8QAILd/lN1qpUYN9WpbP6b6eiu/xIgGFXWaztB
/ygHEZ2Ve/W3YgwAEHnBiVbe18HEiAApi5LKNbU+39oOEfwWANjG2WdqjM9M2Xo/O/FlhbgHrJVS
TuvW69UcWyjwyA0flrwgzbSFpETH+VoSWjfcgtpm39Fjd0Q0HTlVC71LQ/6J06CYBLz9YA08wtPb
sy9Zx2Shi3tQZZyOS1AnD6NPw4Iwmya2JLb5GWYh2XFDmMUSBZda6kDmcDp9e8cYzcWRDI4eLmGA
g+tmnEvzG98qajowNRrW67VjGNkgaqXT924Y6R80eFBJE5usksrLyW/uNGN6XjOzcncLnqTF4rIp
D9u3k57GwnqmIJjzsOylPx6upexZXW35m/sRLmgMjKDJM5Q17jTnky41ic8L5TK4pdf3Q31KvvpW
sTZalgIBEqEeUc/8TwFbLZJ6D5mfxeUEeUMuoKAsXGav/9TGR7TFK0KEgP1OsRWlMbIgSv4o4n9Q
yO+0OCZGspWIk+2GjpE3pSO/7mPq/BTKsS9z9I+RBHJQdf5Lemhho/fXQDj17ILh3vE+23W3lk0k
bNkNF8tEqexdQXzPw/Lgmz6kWAOWw9l4ApR+HvPTKx6ASKZbmCU6kro/kT335qDbdBoB6Opt7EMz
ibF2mZ76/ZSwuBO0OtPgqydEieCQamfHvZKzxsPiEHGwXMVIeau36ohpSgVktWmHP5diElupxasg
8pfjNTUzkPts+geY8rjKqD+XdFhPAZaeCF4D8Q9cRTrdF6h9CRWeo4vlrztDq9Z/AQrxGLcODPk7
e4Ap2A5kkCU+gbQLEYQYSuxgjlYFeeFC1fbD9MYXq2xnpHpZ0pVoWJs6SyhqJTDlOKcg8pVs7HSn
EYh3PFc3U3V1Q9DpiJGg2HZgO4LcHJexhfKSIPPzS1mvDSgsHqDM30FKW3Ho733AiSy6VTH31oM0
dHXf00rJKkujZsDdWZ6ESqgCZD+yh4u1blvbvYxAWCpOTxcY3Wc7yyy8Z9nOG43t2/nI4QnrLTkE
bHdeAKcKYpwPZWMDkaRsBfv6fIvoc0lpiRYXvp/dTvw2OcGT1EekVOktGE7Q4+xHTi1lEPy0jKoP
zgIXfBh5D/yxRhVQCz9wlmpkemC7BEgXJgS09f6fXQCX7Uy/lhEr29704Vcml8fZhtO5bO2uvQ2o
NxZ8k2ZttvwcQZ4Ekb7AfpLFMFNbW6fC1stp6CWLxGSdAlh6Se2+u7ZmBbEE32in+vZXTVlmpQl9
/5hsujej+5Kd0/8ctl8vbXO2ro+63RylhAdR8NCKkyYJilBp35bVIgQRJlZckNW5cL1+VYjVFynh
GC7HYn2UylICMhtUkKYV9nobYzh8R5NHS66fP/ketuezHIx+AWfQbVam3xtamujl3MCh9Pc4gdi9
0DS6QH9xa3HSKMdSF3VL889t6I1ZsW0oP1MEMMu0hBYg239YPrZI0ZRVRXEdImMeRp05uZ7NJQNK
OKbSKQes/UsaakVFoT15gCF5eI9gEhsAwLbIhdVEJuHCO39nEk6RCJMZokebUofuKPzTcX5m4Cqs
JwA5B+caKh1iU0Xqf+Rosb0CXskbqWwiV3bK+n2Tdjovvyh1JrMwoCjm6V9tTG5umDV6NLmE9GUG
OVEddkdTu6NBgVqRFOGYuEngF6UXnVcddwPEVx0o05f2RwuWcIMDxXB9zHIeyMGwV7n5rTDjdJWJ
ksuTcqVody0/MajmmBwLQs4jC7HmQDOgaa4iBaI3zJiq3LROEyczSKQ3NNwHciKbb2T6AG7YRMNv
CxDC1+zGWWBTPhZUskmXntGStYIxZweLi+AGdHpLLbm/ItJjeVieYbhbvWJhRhimUUGC+owEXSmf
Ovbhoju0tYdiZkigTvwwEeYdqcazMrRLobzqJElQngrJJZvSEKQm4EwzM65ck+KHDBuAQ55mZIoX
ZVj0zuE3OaaTxnjP4DKwv8PRdLhFtyx+CJhNqCfjwhe60gMkkvFQM3ZKuKMaS/UNExOFAKhsW0n1
l7fyOeMEs5xRAXXrr8CUc5m3MxopEpEZjfdQL1IcZTQENw5wvQbqGD82Rhh3mwkTbpGGaiPhN+5u
q5xVLcC4AQA22so7pSUN9Q6D6BsYdT+iDbY9Rcd2dEZq4+d92h/E7RYeHB8ynal2eHF7U1U7d/av
IT/FhU4vZehtIc0sy6/KRQGY3lypf71vTdyuxgmSJIMOqUgeq11nKVEdEKnYdUrvWPX8fvHq+B1D
MLfCrDmyAQvPDV2D2dfKKfSuoQfbL2UIrFRvaq3t+3v7RSmBiShYwzVVSALCcECTgxQ3O1Rs5Dj3
L7aeL+xbskwar6bagzMK2nCbGOmSaRn6VpPvDeDRm9oeZzO29UCm72nDpP8NFDvlO/LaxRP4eKjV
ljDVQYVYXYKNbjkDRnjDPN3y6zHnSjV0gsmmrVenGwG/6k3z93neudFtVAOG2NOAUCIXn1wR6EH5
BbHIB2m8erxE0MS+EKIHjHbEu3flrB4rIlOddv7SDaubHpt9e0hXf2SFFdLDz7WMRaeNiMTvP3Pc
9Geb+wvJOHu3O5XZ4vDN86URBIf2DunGMZSlju8UKciZt94KxDaAn6+cRXJqvhKm/gJnU8N8At9X
axnl4oh6IFu+cEfUytH3ziH7CnFn1hjO0WwRGVi8lkfHXl6tTi+mWqQ2cWuOcxNpY3GYTZwW4SOy
GDnkafr7vW3xe2Atq0NYgY5UizLKK87iusmnhG7rMtHDxmGF79eewGXIQyZG8K25fBbjjzVx+dMa
t2TQ1N7SM08rDsItNzOdM5IKl7MR55ZJcdizoKkZ8s7wmJfs2RqX0JxGDqaqbZ5B3LLVoOhsOzyd
15qomCrSmATacWihGA8ZQcl4UMHzV3X4MTxUsCo7+tT38XvQ0erh/uzhVY+E1dcBilnSwt6Ntl19
yIzqLb09X8Rs6KxhocS+pYmMzcRpEFm0iPIosOLT/bfq8aPyqRZxbZ85PDPq19e/qZNQIMv0dSKm
djz7Gn04Rd2DwkwtXhA3QeGwTZpajwfb8jJTFhoQ9jhYw3ovUlF+lohS7x3cElVDYJS/sflP048r
8u2Sx8L8DpxRYSMY5IbXKXnCMUECmwUkjznhF5DTLL4RImOHPLGXb4rCx3BZR2rhrOWKOE9lOZuK
Dg1ADrts6OLGCbjlazM7fdK34SMdvJoYyqyR2/YSFjhJrpQ4fhX/QzHwEryaaCLFMcdH0K+zyLB2
3sJhP0MHGCBChUUS1rEzY9H05ehQodatAK7Fa5wS8QIqbABt4i9YYJfkS5Qmn4/raV54aGqZcg9b
bLSdV1PExHRHBtFIB8Nq3Da/IN4H6Z3+aByaBb5pUS7xbVd7giPLl+4u+KxYVhei0pZXPVc8QDQx
JrhYu4E4EwS/EMf8ss4IpQoqwX+c2lnFIeAOgghks/pvZc5mDJcUAMSryoZzwCQG9EIxc4MIJkdx
Ir0PsBmFgG//w2//HaTxJc3MHs80I3K/zJgtSmKEWPLcXmKgMtIznXCFW4FSHQIMH9vMfcSzSSlk
Pic6RmpGtFzG1jqfCvtO5l1Ppw94/R8zB2caO9OF046OgWDsSt0cCtPaowydGcwfu5Vv8JoYXsiy
fNR/QeXeinyR9vppkDDJCTIcy5X64A9GQcd9Gb0MXwkOdl/6vvNpx3lg1l86D1CSeylJXfjftyFQ
GuM+e4qcXRALTPgvx79v4GHvxASAC6oNDyY0S3nhza3kLAQGoGdGv5qDcqHoki768bt6aTb6Pjwt
6P+yfwcDSB8emw==
`protect end_protected
